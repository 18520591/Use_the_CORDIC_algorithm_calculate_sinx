module Ram(Out, i, clk, reset);
	input [7:0] i;
	input clk, reset;
	output [31:0] Out;
	
	reg [31:0] arctan [0:21];
	always @ (posedge clk, posedge reset)
	begin
		if(reset)
		begin
			arctan[0] <= 32'b01000010001101000000000000000000;
			arctan[1] <= 32'b01000001110101001000010100111001;
			arctan[2] <= 32'b01000001011000001001010001110100;
			arctan[3] <= 32'b01000000111001000000000000100010;
			arctan[4] <= 32'b01000000011001001110001010101001;
			arctan[5] <= 32'b00111111111001010001101111001010;
			arctan[6] <= 32'b00111111011001010010101000011010;
			arctan[7] <= 32'b00111110111001010010110110101111;
			arctan[8] <= 32'b00111110011001010010111010010100;
			arctan[9] <= 32'b00111101111001010010111011001101;
			arctan[10] <= 32'b00111101011001010010111011011100;
			arctan[11] <= 32'b00111100111001010010111011011111;
			arctan[12] <= 32'b00111100011001010010111011100000;
			arctan[13] <= 32'b00111011111001010010111011100000;
			arctan[14] <= 32'b00111011011001010010111011100000;
			arctan[15] <= 32'b00111011111101010100011100011101;
			arctan[16] <= 32'b00111010011001010010111011100000;
			arctan[17] <= 32'b00111001111001010010111011100000;
			arctan[18] <= 32'b00111001011001010010111011100000;
			arctan[19] <= 32'b00111000111001010010111011100000;
			arctan[20] <= 32'b00111000011001010010111011100000;
		end
	end
	assign Out = arctan[i];
endmodule